module TD4 (
    input CLK,
    input CLR,

    input [7:0] D,
    output [3:0] A
);
    
endmodule
